library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library wave;
use wave.wave_array_pkg.all;

library osc;


entity noise_source is 
    port (
        clk                     : in  std_logic;
        reset                   : in  std_logic;
        config                  : in  t_config;
        next_sample             : in  std_logic;
        output_samples          : out t_mono_sample_array(POLYPHONY_MAX - 1 downto 0)
    );
end entity;


architecture arch of noise_source is

    -- Magic numbers.
    constant SHIFT_IN   : integer := 6; -- Right shift input samples to brown noise accumulator by this amount
    constant SHIFT_LEAK : integer := 10; -- Decrease sum by this frac each cycle to avoid overflow. 

    type t_state is (idle, sample_bits, finalize_0, finalize_1);

    type t_noise_reg is record
        state                   : t_state;
        bit_count               : integer range 0 to SAMPLE_SIZE - 1;
        voice_count             : integer range 0 to POLYPHONY_MAX - 1;
        output_samples          : t_mono_sample_array(POLYPHONY_MAX - 1 downto 0);
        sample_buffers          : t_mono_sample_array(POLYPHONY_MAX - 1 downto 0);
        noise_select            : std_logic;
        sum                     : t_mono_sample;
    end record;

    constant REG_INIT : t_noise_reg := (
        state                   => idle,
        bit_count               => 0,
        voice_count             => 0,
        output_samples          => (others => (others => '0')),
        sample_buffers          => (others => (others => '0')),
        noise_select            => '0',
        sum                     => (others => '0')
    );

    signal r, r_in              : t_noise_reg;
    signal s_read_enable        : std_logic;
    signal s_output_valid       : std_logic;
    signal s_output_data        : std_logic;    

begin

    lfsr : entity osc.lfsr32 
    port map (
        clk                     => clk,
        reset                   => reset,
        read_enable             => s_read_enable,
        output_valid            => s_output_valid,
        output_data             => s_output_data
    );


    comb_process : process (r, config, next_sample, s_output_valid, s_output_data)
    begin

        r_in <= r;
        r_in.noise_select <= config.noise_select;
        s_read_enable <= '0';

        output_samples <= r.output_samples;
        
        if r.state = idle then
            if next_sample = '1' then 
                r_in.output_samples <= r.sample_buffers;
                r_in.bit_count <= 0;                    
                r_in.voice_count <= 0;
                s_read_enable <= '1';
                r_in.state <= sample_bits;
            end if;
           
        elsif r.state = sample_bits then 

            if s_output_valid = '1' then 

                r_in.sample_buffers(r.voice_count)(r.bit_count) <= s_output_data;
                
                if r.bit_count < SAMPLE_SIZE - 1 then 
                    s_read_enable <= '1';
                    r_in.bit_count <= r.bit_count + 1;
                else 
                    r_in.state <= finalize_0;
                end if;
            end if;

        elsif r.state = finalize_0 then

            r_in.bit_count <= 0;

            -- Brown noise is generated by integrating the (shifted) noise samples. 
            if r.noise_select = '0' then

                r_in.sum <= r.output_samples(r.voice_count) + shift_right(r.sample_buffers(r.voice_count), SHIFT_IN);

            -- White noise is just the samples directly. 
            -- But divided by two to make the amplitude similar to the brown noise.
            else 
                r_in.sum <= r.sample_buffers(r.voice_count);
            end if;

            r_in.state <= finalize_1;

        elsif r.state = finalize_1 then

            r_in.sample_buffers(r.voice_count) <= r.sum - shift_right(r.sum, SHIFT_LEAK);

            if r.voice_count < POLYPHONY_MAX - 1 then 
                r_in.voice_count <= r.voice_count + 1;
                s_read_enable <= '1';
                r_in.state <= sample_bits;
            else 
                r_in.state <= idle;
            end if;
        end if;

    end process;


    reg_process : process (clk)
    begin
        if rising_edge(clk) then
            if reset = '1' then
                r <= REG_INIT;
            else
                r <= r_in;
            end if;
        end if;
    end process;

end architecture;
